// megafunction wizard: %Test-Pattern Generator v13.0%
// GENERATION: XML
// test_pattern_gen_ip.v

// Generated using ACDS version 13.0sp1 232 at 2023.01.28.15:21:26

`timescale 1 ps / 1 ps
module test_pattern_gen_ip (
		input  wire        clk,           //             clock_reset.clk
		input  wire        reset,         //       clock_reset_reset.reset
		input  wire        ready,         // avalon_generator_source.ready
		output wire [23:0] data,          //                        .data
		output wire        startofpacket, //                        .startofpacket
		output wire        endofpacket,   //                        .endofpacket
		output wire        valid          //                        .valid
	);

	test_pattern_gen_ip_0002 test_pattern_gen_ip_inst (
		.clk           (clk),           //             clock_reset.clk
		.reset         (reset),         //       clock_reset_reset.reset
		.ready         (ready),         // avalon_generator_source.ready
		.data          (data),          //                        .data
		.startofpacket (startofpacket), //                        .startofpacket
		.endofpacket   (endofpacket),   //                        .endofpacket
		.valid         (valid)          //                        .valid
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2023 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_up_avalon_video_test_pattern" version="13.0" >
// Retrieval info: 	<generic name="width" value="720" />
// Retrieval info: 	<generic name="height" value="720" />
// Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone II" />
// Retrieval info: </instance>
// IPFS_FILES : test_pattern_gen_ip.vo
// RELATED_FILES: test_pattern_gen_ip.v, test_pattern_gen_ip_0002.v
