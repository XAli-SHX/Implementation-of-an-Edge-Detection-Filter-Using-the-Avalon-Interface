library verilog;
use verilog.vl_types.all;
entity CounterDualPort_tb is
end CounterDualPort_tb;
