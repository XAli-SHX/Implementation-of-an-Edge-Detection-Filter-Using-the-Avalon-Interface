library verilog;
use verilog.vl_types.all;
entity Sobel_AvalonStreaming_tb is
end Sobel_AvalonStreaming_tb;
