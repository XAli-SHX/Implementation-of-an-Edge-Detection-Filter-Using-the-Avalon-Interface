library verilog;
use verilog.vl_types.all;
entity SobelFilter_tb is
end SobelFilter_tb;
