// megafunction wizard: %VGA Controller v13.0%
// GENERATION: XML
// vga_controller_ip.v

// Generated using ACDS version 13.0sp1 232 at 2023.01.28.15:33:47

`timescale 1 ps / 1 ps
module vga_controller_ip (
		input  wire        clk,           //        clock_reset.clk
		input  wire        reset,         //  clock_reset_reset.reset
		input  wire [29:0] data,          //    avalon_vga_sink.data
		input  wire        startofpacket, //                   .startofpacket
		input  wire        endofpacket,   //                   .endofpacket
		input  wire        valid,         //                   .valid
		output wire        ready,         //                   .ready
		output wire        VGA_CLK,       // external_interface.export
		output wire        VGA_HS,        //                   .export
		output wire        VGA_VS,        //                   .export
		output wire        VGA_BLANK,     //                   .export
		output wire        VGA_SYNC,      //                   .export
		output wire [9:0]  VGA_R,         //                   .export
		output wire [9:0]  VGA_G,         //                   .export
		output wire [9:0]  VGA_B          //                   .export
	);

	vga_controller_ip_0002 vga_controller_ip_inst (
		.clk           (clk),           //        clock_reset.clk
		.reset         (reset),         //  clock_reset_reset.reset
		.data          (data),          //    avalon_vga_sink.data
		.startofpacket (startofpacket), //                   .startofpacket
		.endofpacket   (endofpacket),   //                   .endofpacket
		.valid         (valid),         //                   .valid
		.ready         (ready),         //                   .ready
		.VGA_CLK       (VGA_CLK),       // external_interface.export
		.VGA_HS        (VGA_HS),        //                   .export
		.VGA_VS        (VGA_VS),        //                   .export
		.VGA_BLANK     (VGA_BLANK),     //                   .export
		.VGA_SYNC      (VGA_SYNC),      //                   .export
		.VGA_R         (VGA_R),         //                   .export
		.VGA_G         (VGA_G),         //                   .export
		.VGA_B         (VGA_B)          //                   .export
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2023 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_up_avalon_video_vga_controller" version="13.0" >
// Retrieval info: 	<generic name="board" value="DE2" />
// Retrieval info: 	<generic name="device" value="VGA Connector" />
// Retrieval info: 	<generic name="underflow_flag" value="false" />
// Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone II" />
// Retrieval info: </instance>
// IPFS_FILES : vga_controller_ip.vo
// RELATED_FILES: vga_controller_ip.v, altera_up_avalon_video_vga_timing.v, vga_controller_ip_0002.v
