// megafunction wizard: %Character Buffer for VGA Display v13.0%
// GENERATION: XML
// vga_display_cb_ip.v

// Generated using ACDS version 13.0sp1 232 at 2023.01.28.15:32:05

`timescale 1 ps / 1 ps
module vga_display_cb_ip (
		input  wire        clk,                  //               clock_reset.clk
		input  wire        reset,                //         clock_reset_reset.reset
		input  wire        ctrl_address,         // avalon_char_control_slave.address
		input  wire [3:0]  ctrl_byteenable,      //                          .byteenable
		input  wire        ctrl_chipselect,      //                          .chipselect
		input  wire        ctrl_read,            //                          .read
		input  wire        ctrl_write,           //                          .write
		input  wire [31:0] ctrl_writedata,       //                          .writedata
		output wire [31:0] ctrl_readdata,        //                          .readdata
		input  wire        buf_byteenable,       //  avalon_char_buffer_slave.byteenable
		input  wire        buf_chipselect,       //                          .chipselect
		input  wire        buf_read,             //                          .read
		input  wire        buf_write,            //                          .write
		input  wire [7:0]  buf_writedata,        //                          .writedata
		output wire [7:0]  buf_readdata,         //                          .readdata
		output wire        buf_waitrequest,      //                          .waitrequest
		input  wire [12:0] buf_address,          //                          .address
		input  wire        stream_ready,         //        avalon_char_source.ready
		output wire        stream_startofpacket, //                          .startofpacket
		output wire        stream_endofpacket,   //                          .endofpacket
		output wire        stream_valid,         //                          .valid
		output wire [29:0] stream_data           //                          .data
	);

	vga_display_cb_ip_0002 vga_display_cb_ip_inst (
		.clk                  (clk),                  //               clock_reset.clk
		.reset                (reset),                //         clock_reset_reset.reset
		.ctrl_address         (ctrl_address),         // avalon_char_control_slave.address
		.ctrl_byteenable      (ctrl_byteenable),      //                          .byteenable
		.ctrl_chipselect      (ctrl_chipselect),      //                          .chipselect
		.ctrl_read            (ctrl_read),            //                          .read
		.ctrl_write           (ctrl_write),           //                          .write
		.ctrl_writedata       (ctrl_writedata),       //                          .writedata
		.ctrl_readdata        (ctrl_readdata),        //                          .readdata
		.buf_byteenable       (buf_byteenable),       //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (buf_chipselect),       //                          .chipselect
		.buf_read             (buf_read),             //                          .read
		.buf_write            (buf_write),            //                          .write
		.buf_writedata        (buf_writedata),        //                          .writedata
		.buf_readdata         (buf_readdata),         //                          .readdata
		.buf_waitrequest      (buf_waitrequest),      //                          .waitrequest
		.buf_address          (buf_address),          //                          .address
		.stream_ready         (stream_ready),         //        avalon_char_source.ready
		.stream_startofpacket (stream_startofpacket), //                          .startofpacket
		.stream_endofpacket   (stream_endofpacket),   //                          .endofpacket
		.stream_valid         (stream_valid),         //                          .valid
		.stream_data          (stream_data)           //                          .data
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2023 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_up_avalon_video_character_buffer_with_dma" version="13.0" >
// Retrieval info: 	<generic name="vga_device" value="On-board VGA DAC" />
// Retrieval info: 	<generic name="enable_transparency" value="false" />
// Retrieval info: 	<generic name="color_bits" value="1-bit" />
// Retrieval info: 	<generic name="resolution" value="80 x 60" />
// Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone II" />
// Retrieval info: </instance>
// IPFS_FILES : vga_display_cb_ip.vo
// RELATED_FILES: vga_display_cb_ip.v, altera_up_video_128_character_rom.v, altera_up_video_fb_color_rom.v, vga_display_cb_ip_0002.v
