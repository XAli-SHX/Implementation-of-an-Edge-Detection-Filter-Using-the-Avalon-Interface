library verilog;
use verilog.vl_types.all;
entity EdgeDetector_tb is
end EdgeDetector_tb;
