// megafunction wizard: %Edge Detection v13.0%
// GENERATION: XML
// edge_detector_ip.v

// Generated using ACDS version 13.0sp1 232 at 2023.01.28.15:20:01

`timescale 1 ps / 1 ps
module edge_detector_ip (
		input  wire       clk,               //                  clock_reset.clk
		input  wire       reset,             //            clock_reset_reset.reset
		input  wire [7:0] in_data,           //   avalon_edge_detection_sink.data
		input  wire       in_startofpacket,  //                             .startofpacket
		input  wire       in_endofpacket,    //                             .endofpacket
		input  wire       in_valid,          //                             .valid
		output wire       in_ready,          //                             .ready
		input  wire       out_ready,         // avalon_edge_detection_source.ready
		output wire [7:0] out_data,          //                             .data
		output wire       out_startofpacket, //                             .startofpacket
		output wire       out_endofpacket,   //                             .endofpacket
		output wire       out_valid          //                             .valid
	);

	edge_detector_ip_0002 edge_detector_ip_inst (
		.clk               (clk),               //                  clock_reset.clk
		.reset             (reset),             //            clock_reset_reset.reset
		.in_data           (in_data),           //   avalon_edge_detection_sink.data
		.in_startofpacket  (in_startofpacket),  //                             .startofpacket
		.in_endofpacket    (in_endofpacket),    //                             .endofpacket
		.in_valid          (in_valid),          //                             .valid
		.in_ready          (in_ready),          //                             .ready
		.out_ready         (out_ready),         // avalon_edge_detection_source.ready
		.out_data          (out_data),          //                             .data
		.out_startofpacket (out_startofpacket), //                             .startofpacket
		.out_endofpacket   (out_endofpacket),   //                             .endofpacket
		.out_valid         (out_valid)          //                             .valid
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2023 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_up_avalon_video_edge_detection" version="13.0" >
// Retrieval info: 	<generic name="width" value="720" />
// Retrieval info: 	<generic name="intensity" value="1" />
// Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone II" />
// Retrieval info: </instance>
// IPFS_FILES : edge_detector_ip.vo
// RELATED_FILES: edge_detector_ip.v, altera_up_edge_detection_gaussian_smoothing_filter.v, altera_up_edge_detection_sobel_operator.v, altera_up_edge_detection_nonmaximum_suppression.v, altera_up_edge_detection_hysteresis.v, altera_up_edge_detection_pixel_info_shift_register.v, altera_up_edge_detection_data_shift_register.v, edge_detector_ip_0002.v
