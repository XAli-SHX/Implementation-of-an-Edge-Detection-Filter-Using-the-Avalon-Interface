library verilog;
use verilog.vl_types.all;
entity Rgb2Gray_tb is
end Rgb2Gray_tb;
