library verilog;
use verilog.vl_types.all;
entity AnyImage_tb is
end AnyImage_tb;
